class Baseinstr ;//extends uvm_object;
static reg[31:0] instr;

endclass
